`timescale 1ns / 1ps

module ROM(ROM_address,
			  ROM_data
    );

input [7:0] ROM_address;
output [7:0] ROM_data;

	reg [7:0] Cel [255:0];

		initial begin
	
		Cel[0] = 8'b00000000;
// Calculate Image Full Size
Cel[1] = 8'b00000001;
Cel[2] = 8'b00000000;
Cel[3] = 8'b00001101;
Cel[4] = 8'b10010001;
Cel[5] = 8'b00000100;
Cel[6] = 8'b00000001;
Cel[7] = 8'b00000000;
Cel[8] = 8'b00001110;
Cel[9] = 8'b00001101;
Cel[10] = 8'b00000010;
Cel[11] = 8'b00000000;
Cel[12] = 8'b00000000;
//Image Processing Start
Cel[13] = 8'b00000001;
Cel[14] = 8'b00000000;
Cel[15] = 8'b00000011;
Cel[16] = 8'b00000010;
Cel[17] = 8'b00000000;
Cel[18] = 8'b00000100;
Cel[19] = 8'b00000010;
Cel[20] = 8'b00000000;
Cel[21] = 8'b00000101;
Cel[22] = 8'b00000001;
Cel[23] = 8'b00000000;
Cel[24] = 8'b00001001;
Cel[25] = 8'b00000100;
Cel[26] = 8'b00000001;
Cel[27] = 8'b00000000;
Cel[28] = 8'b00000010;
Cel[29] = 8'b00000101;
Cel[30] = 8'b00000001;
Cel[31] = 8'b00000000;
Cel[32] = 8'b00000011;
Cel[33] = 8'b00001111;
Cel[34] = 8'b00001110;
Cel[35] = 8'b00000010;
Cel[36] = 8'b00000000;
Cel[37] = 8'b00000110;
Cel[38] = 8'b00000001;
Cel[39] = 8'b00000000;
Cel[40] = 8'b00000000;
Cel[41] = 8'b00000100;
Cel[42] = 8'b00000001;
Cel[43] = 8'b00000000;
Cel[44] = 8'b00000011;
Cel[45] = 8'b00001101;
Cel[46] = 8'b00000010;
Cel[47] = 8'b00000000;
Cel[48] = 8'b00000111;
Cel[49] = 8'b00000001;
Cel[50] = 8'b00000000;
Cel[51] = 8'b00000001;
Cel[52] = 8'b00000100;
Cel[53] = 8'b00000001;
Cel[54] = 8'b00000000;
Cel[55] = 8'b00000111;
Cel[56] = 8'b00001110;
Cel[57] = 8'b00001110;
Cel[58] = 8'b00000010;
Cel[59] = 8'b00000000;
Cel[60] = 8'b00001000;

//Start Of First Loop

Cel[61] = 8'b00001000;
Cel[62] = 8'b00000000;
Cel[63] = 8'b00000101;
Cel[64] = 8'b00001010;
Cel[65] = 8'b00000100;
Cel[66] = 8'b00000001;
Cel[67] = 8'b00000000;
Cel[68] = 8'b00000101;
Cel[69] = 8'b00001100;
Cel[70] = 8'b00000010;
Cel[71] = 8'b00000000;
Cel[72] = 8'b00000101;
Cel[73] = 8'b00001000;
Cel[74] = 8'b00000000;
Cel[75] = 8'b00000101;
Cel[76] = 8'b00001011;
Cel[77] = 8'b00001101;
Cel[78] = 8'b00000100;
Cel[79] = 8'b00000001;
Cel[80] = 8'b00000000;
Cel[81] = 8'b00000101;
Cel[82] = 8'b00001100;
Cel[83] = 8'b00000010;
Cel[84] = 8'b00000000;
Cel[85] = 8'b00000101;
Cel[86] = 8'b00001000;
Cel[87] = 8'b00000000;
Cel[88] = 8'b00000101;
Cel[89] = 8'b00001010;
Cel[90] = 8'b00001101;
Cel[91] = 8'b00001001;
Cel[92] = 8'b00000000;
Cel[93] = 8'b00000100;
Cel[94] = 8'b00000001;
Cel[95] = 8'b00000000;
Cel[96] = 8'b00000100;
Cel[97] = 8'b00001100;
Cel[98] = 8'b00000010;
Cel[99] = 8'b00000000;
Cel[100] = 8'b00000100;
Cel[101] = 8'b00000010;
Cel[102] = 8'b00000000;
Cel[103] = 8'b00000101;
Cel[104] = 8'b00000100;
Cel[105] = 8'b00000001;
Cel[106] = 8'b00000000;
Cel[107] = 8'b00000110;
Cel[108] = 8'b00001110;
Cel[109] = 8'b00000111;
Cel[110] = 8'b00111101;
//ROW wise
Cel[111] = 8'b00000001;
Cel[112] = 8'b00000000;
Cel[113] = 8'b00000110;
Cel[114] = 8'b00001111;
Cel[115] = 8'b00000010;
Cel[116] = 8'b00000000;
Cel[117] = 8'b00000110;
Cel[118] = 8'b00000001;
Cel[119] = 8'b00000000;
Cel[120] = 8'b00000100;
Cel[121] = 8'b00001100;
Cel[122] = 8'b00001100;
Cel[123] = 8'b00000010;
Cel[124] = 8'b00000000;
Cel[125] = 8'b00000100;
Cel[126] = 8'b00000010;
Cel[127] = 8'b00000000;
Cel[128] = 8'b00000101;
Cel[129] = 8'b00000100;
Cel[130] = 8'b00000001;
Cel[131] = 8'b00000000;
Cel[132] = 8'b00000111;
Cel[133] = 8'b00001110;
Cel[134] = 8'b00000111;
Cel[135] = 8'b00111101;
/*************END of LOOP_1*******************************/
Cel[136] = 8'b00000001;
Cel[137] = 8'b00000000;
Cel[138] = 8'b00000011;
Cel[139] = 8'b00000010;
Cel[140] = 8'b00000000;
Cel[141] = 8'b00000100;
Cel[142] = 8'b00000010;
Cel[143] = 8'b00000000;
Cel[144] = 8'b00000101;
Cel[145] = 8'b00000001;
Cel[146] = 8'b00000000;
Cel[147] = 8'b00001001;
Cel[148] = 8'b00000100;
Cel[149] = 8'b00000001;
Cel[150] = 8'b00000000;
Cel[151] = 8'b00000010;
Cel[152] = 8'b00000101;
Cel[153] = 8'b00000001;
Cel[154] = 8'b00000000;
Cel[155] = 8'b00000011;
Cel[156] = 8'b00001111;
Cel[157] = 8'b00001110;
Cel[158] = 8'b00000010;
Cel[159] = 8'b00000000;
Cel[160] = 8'b00000110;
/**********Start of LOOP_2******************/
Cel[161] = 8'b00001000;
Cel[162] = 8'b00000000;
Cel[163] = 8'b00000101;
Cel[164] = 8'b00001010;
Cel[165] = 8'b00000100;
Cel[166] = 8'b00000001;
Cel[167] = 8'b00000000;
Cel[168] = 8'b00000101;
Cel[169] = 8'b00001111;
Cel[170] = 8'b00000010;
Cel[171] = 8'b00000000;
Cel[172] = 8'b00000101;
Cel[173] = 8'b00001000;
Cel[174] = 8'b00000000;
Cel[175] = 8'b00000101;
Cel[176] = 8'b00001011;
Cel[177] = 8'b00001101;
Cel[178] = 8'b00000100;
Cel[179] = 8'b00000001;
Cel[180] = 8'b00000000;
Cel[181] = 8'b00000101;
Cel[182] = 8'b00001111;
Cel[183] = 8'b00000010;
Cel[184] = 8'b00000000;
Cel[185] = 8'b00000101;
Cel[186] = 8'b00001000;
Cel[187] = 8'b00000000;
Cel[188] = 8'b00000101;
Cel[189] = 8'b00001010;
Cel[190] = 8'b00001101;
Cel[191] = 8'b00001001;
Cel[192] = 8'b00000000;
Cel[193] = 8'b00000100;
Cel[194] = 8'b00000001;
Cel[195] = 8'b00000000;
Cel[196] = 8'b00000100;
Cel[197] = 8'b00001100;
Cel[198] = 8'b00000010;
Cel[199] = 8'b00000000;
Cel[200] = 8'b00000100;
Cel[201] = 8'b00000010;
Cel[202] = 8'b00000000;
Cel[203] = 8'b00000101;
Cel[204] = 8'b00000100;
Cel[205] = 8'b00000001;
Cel[206] = 8'b00000000;
Cel[207] = 8'b00001000;
Cel[208] = 8'b00001110;
Cel[209] = 8'b00000111;
Cel[210] = 8'b10100001;
// Store Image Start Here
Cel[211] = 8'b00000001;
Cel[212] = 8'b00000000;
Cel[213] = 8'b00000111;
Cel[214] = 8'b00001111;
Cel[215] = 8'b00000010;
Cel[216] = 8'b00000000;
Cel[217] = 8'b00001010;
Cel[218] = 8'b00000010;
Cel[219] = 8'b00000000;
Cel[220] = 8'b00001011;
Cel[221] = 8'b00000001;
Cel[222] = 8'b00000000;
Cel[223] = 8'b00000011;
Cel[224] = 8'b00000010;
Cel[225] = 8'b00000000;
Cel[226] = 8'b00000100;
Cel[227] = 8'b00000010;
Cel[228] = 8'b00000000;
Cel[229] = 8'b00000101;
Cel[230] = 8'b00000001;
Cel[231] = 8'b00000000;
Cel[232] = 8'b00001001;
Cel[233] = 8'b00001011;
Cel[234] = 8'b00000100;
Cel[235] = 8'b00000001;
Cel[236] = 8'b00000000;
Cel[237] = 8'b00000011;
Cel[238] = 8'b00001111;
Cel[239] = 8'b00001110;
Cel[240] = 8'b00000010;
Cel[241] = 8'b00000000;
Cel[242] = 8'b00000110;
		//End of Process
		Cel[243] = 8'b10101010;

	end
	
assign ROM_data =Cel[ROM_address];

endmodule
