`timescale 1ns / 1ps
module ControlUnit(Z_EN,RAM_en,REG_INC,Z,MPC,clk,Addr,JMPC,ALU,C,B,M,End_of_process
    );

	input clk,Z;
	input [7:0] MPC;
	
	output [7:0] Addr;
	output [3:0] ALU;
	output [5:0] C;
	output [2:0] B;
	output [1:0] M;
	output [2:0] REG_INC;
	output JMPC;
	output RAM_en;
	output Z_EN;
	output End_of_process;
	
	reg End_of_process;
	reg [28:0] CL_MEM [511:0];
	reg [28:0] MIR;
	//Instructions
	
//-------------------------------------------------------
	initial 
	begin
	
	MIR = 29'b0_0_00000000_000000_000_000_0000_000;

	//assign {JMPC,Z_EN,Addr,C,REG_INC,B,ALU,RAM_en,M} = MIR; 
			/*3'b000 : B_bus <= B_bus;
			3'b001 : B_bus <= GP;
			3'b010 : B_bus <= PC;
			3'b011 : B_bus <= GP2;
			3'b100 : B_bus <= MDR;
			3'b101 : B_bus <= MAR;
			3'b110 : B_bus <= IR;
			3'b111 : B_bus <=  16'bz;*/
	//1.Nop
	 CL_MEM[9'b000000000]= 29'b1_0_00000000_000000_001_000_0000_000;	
	 
	 //2.Load AC from Memory (AC <- M[T] -0000 0001 T1,T2)
	 CL_MEM[9'b000000001]= 29'b0_0_00010001_000000_001_000_0000_000;
	 CL_MEM[9'b00001_0001]= 29'b0_0_00010010_000001_001_110_1011_000;
	 CL_MEM[9'b000010010]= 29'b0_0_00010011_010000_000_110_0100_000;
	 CL_MEM[9'b000010011]= 29'b0_0_00010100_000000_000_000_0000_000;
	 CL_MEM[9'b000010100]= 29'b0_0_00010101_000000_000_000_0000_101;
	 CL_MEM[9'b000010101]= 29'b0_0_00010111_000000_000_000_0000_101;
	 CL_MEM[9'b000010111]= 29'b0_0_00000000_000001_000_100_0011_000;
		
	 //3.LOAD Memory with AC (M[T] <- AC -0000 0010 T1,T2)
	 CL_MEM[9'b000000010]= 29'b0_0_00100000_001000_000_000_0010_000;
	 CL_MEM[9'b00010_0000]= 29'b0_0_00100001_000000_001_000_0000_000;
	 CL_MEM[9'b000100001]= 29'b0_0_00100010_000001_001_110_1011_000;
	 CL_MEM[9'b000100010]= 29'b0_0_00100011_010000_000_110_0100_000;
	 CL_MEM[9'b000100011]= 29'b0_0_00100100_000000_000_000_0000_110;
	 CL_MEM[9'b000100100]= 29'b0_0_00100101_000000_000_000_0000_110;
	 CL_MEM[9'b000100101]= 29'b0_0_00000000_000001_000_100_0011_000;
	 
	 
	 //4.Clear AC
	 CL_MEM[9'b000000011]= 29'b0_0_00000000_000001_000_000_0001_000;
	 
	 //5.MOVE AC GP1
	CL_MEM[9'b000000100]= 29'b0_0_00110000_000010_000_000_0010_000;
	CL_MEM[9'b00011_0000]= 29'b0_0_00000000_000000_000_000_0000_000;
	
	
	 //6.MOVE AC GP1
	CL_MEM[9'b000000101]= 29'b0_0_01000000_100000_000_000_0010_000;
	CL_MEM[9'b00100_0000]= 29'b0_0_00000000_000000_000_000_0000_000;

	//7. JUMPZ
	CL_MEM[9'b000000110]= 29'b0_1_01010000_000000_000_110_0011_000;
		//If AC = 0;
	CL_MEM[9'b10101_0000]= 29'b0_1_01010001_000100_000_110_0011_000;
	CL_MEM[9'b101010001]= 29'b1_0_00000000_000000_001_000_0000_000;
		//If AC != 0;
	CL_MEM[9'b001010000]= 29'b0_0_00000000_000000_001_110_0011_000;
	
	//8. JUMNZ
	CL_MEM[9'b000000111]= 29'b0_1_01100000_000000_000_110_0011_000;
		//If AC != 0;
	CL_MEM[9'b00110_0000]= 29'b0_1_01100001_000100_000_110_0011_000;
	CL_MEM[9'b001100001]= 29'b1_0_00000000_000000_001_000_0000_000;
		//If AC == 0;
	CL_MEM[9'b101100000]= 29'b0_0_00000000_000000_001_110_0011_000;
	
	//8. Load AC  AC<= M[M[T,T]]
	 CL_MEM[9'b000001000]= 29'b0_0_01110000_000000_001_000_0000_000;
	 CL_MEM[9'b001110000]= 29'b0_0_01110001_000001_001_110_1011_000;
	 CL_MEM[9'b001110001]= 29'b0_0_01110010_010000_000_110_0100_000;
	 CL_MEM[9'b001110010]= 29'b0_0_01110011_000000_000_000_0000_000;
	 CL_MEM[9'b001110011]= 29'b0_0_01110100_000000_000_000_0000_101;
	 CL_MEM[9'b001110100]= 29'b0_0_01110101_000000_000_000_0000_101;
	 CL_MEM[9'b001110101]= 29'b0_0_01110110_010000_000_100_0011_000;
	 CL_MEM[9'b001110110]= 29'b0_0_01110111_000000_000_000_0000_101;
	 CL_MEM[9'b001110111]= 29'b0_0_01111000_000000_000_000_0000_101;
	 CL_MEM[9'b001111000]= 29'b0_0_00000000_000001_000_100_0011_000;

	//9. Store AC - M[M[T,T]] <= AC
	 CL_MEM[9'b000001001]= 29'b0_0_10000000_001000_000_000_0010_000;
	 CL_MEM[9'b010000000]= 29'b0_0_10000001_000000_001_000_0000_000;
	 CL_MEM[9'b010000001]= 29'b0_0_10000010_000001_001_110_1011_000;
	 CL_MEM[9'b010000010]= 29'b0_0_10000011_010000_000_110_0100_000;
	 CL_MEM[9'b010000011]= 29'b0_0_10000100_000001_000_100_0011_000;
	 CL_MEM[9'b010000100]= 29'b0_0_10000101_000000_000_000_0000_101;
	 CL_MEM[9'b010000101]= 29'b0_0_10000110_000000_000_000_0000_101;
	 CL_MEM[9'b010000110]= 29'b0_0_10000111_010000_000_100_0011_000;
	 CL_MEM[9'b010000111]= 29'b0_0_10001000_001000_000_000_0010_000;
	 CL_MEM[9'b010001000]= 29'b0_0_10001001_000000_000_000_0000_110;
	 CL_MEM[9'b010001001]= 29'b0_0_00000000_000000_000_000_0000_110;
	
	
	//10.DIV AC by 4
	 CL_MEM[9'b000001010]= 29'b0_0_10010000_000001_000_000_0110_000;
	 CL_MEM[9'b010010000]= 29'b0_0_00000000_000000_000_000_0000_000;
	 
	//11.DIV AC by 2
	 CL_MEM[9'b000001011]= 29'b0_0_10100000_000001_000_000_0111_000;
	 CL_MEM[9'b010100000]= 29'b0_0_00000000_000000_000_000_0000_000;
	
	//12. INC AC
	 CL_MEM[9'b000001100]= 29'b0_0_10110000_000001_000_000_1010_000;
	 CL_MEM[9'b010110000]= 29'b0_0_00000000_000000_000_000_0000_000;
	 
	 //13. ADD AC + GP1
	 CL_MEM[9'b000001101]= 29'b0_0_11000000_000001_000_001_0100_000;
	 CL_MEM[9'b011000000]= 29'b0_0_00000000_000000_000_000_0000_000;
	 
	 //14. SUB AC - GP1
	 CL_MEM[9'b000001110]= 29'b0_0_11010000_000001_000_001_0101_000;
	 CL_MEM[9'b011010000]= 29'b0_0_00000000_000000_000_000_0000_000;
	 
	 //15. ADD AC + GP2
	 CL_MEM[9'b000001111]= 29'b0_0_11100000_000001_000_011_0100_000;
	 CL_MEM[9'b011100000]= 29'b0_0_00000000_000000_000_000_0000_000;
	 
	 //16.Shift AC by 8
	 CL_MEM[9'b010010001]= 29'b0_0_10010010_000001_000_000_1100_000;
	 CL_MEM[9'b010010010]= 29'b0_0_00000000_000000_000_000_0000_000;
	 
	 
	 End_of_process=1'b0;
	end
//----------------------------------------------------	
	
	always @ (negedge clk) begin
		MIR = CL_MEM[{Z,MPC}];                               //rlease cl sig in posedge
		
		if(MPC == 8'b10101010)
			begin
				End_of_process<= 1'b1;
			end
		else
			begin
				End_of_process<= 1'b0;
			end
	end
	
	
	assign {JMPC,Z_EN,Addr,C,REG_INC,B,ALU,RAM_en,M} = MIR;  
	//0_0_00000000_000000_000_000_0000_000

endmodule
