`timescale 1ns / 1ps
module Test_UART;

	// Inputs
	reg clk;
	reg PC_RAM_ACT;
	reg RAM_PC_ACT;
	reg PROCESS_ACT;

	// Instantiate the Unit Under Test (UUT)
	Top uut (
		.clk(clk), 
		.PC_RAM_ACT(PC_RAM_ACT), 
		.RAM_PC_ACT(RAM_PC_ACT), 
		.PROCESS_ACT(PROCESS_ACT)
	);

	always #5 clk=~clk;
	
	initial begin
		// Initialize Inputs
		clk = 0;
		PC_RAM_ACT = 0;
		RAM_PC_ACT = 0;
		PROCESS_ACT = 0;
		
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
			#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
			#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
			#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
			#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;

		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
			#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
			#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
			#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
			#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
			#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
			#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
			#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
			#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
			#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
			#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
			#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
			#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
			#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
			#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
			#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
			#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
			#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
			#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
			#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
			#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;
		#0.1 RAM_PC_ACT=~RAM_PC_ACT;		
		#100;
        
		// Add stimulus here

	end
      
endmodule

